library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

package cordic_lib is
    type tupla is array(NATURAL range <>) of SIGNED;
end cordic_lib;