library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.my_library.all;
entity delay is
    port (i_in : in  t_punto;
	  clk : in std_logic;
	  o_out : out t_punto);
end delay;
architecture delay_arq of delay is
signal mem : t_punto := ((x=> (others => '0'),y => (others => '0')));
begin
process (clk)
begin
o_out <= mem;
mem <= i_in;
end process;
end delay_arq;